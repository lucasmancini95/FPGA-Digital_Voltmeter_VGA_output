----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.02.2020 17:28:48
-- Design Name: 
-- Module Name: counter_generic_bis_tb - counter_generic_bis_tb_arq
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity counter_generic_bis_tb is
    Port ( d : in STD_LOGIC);
end counter_generic_bis_tb;

architecture counter_generic_bis_tb_arq of counter_generic_bis_tb is

begin


end counter_generic_bis_tb_arq;
